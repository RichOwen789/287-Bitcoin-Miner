module rev256(in,out);
input [255:0]in;
output [255:0]out;
wire [255:0]out;
assign out[0] = in[255];                                                                                                                                                                                                                                
assign out[1] = in[254];                                                                                                                                                                                                                                
assign out[2] = in[253];                                                                                                                                                                                                                                
assign out[3] = in[252];                                                                                                                                                                                                                                
assign out[4] = in[251];                                                                                                                                                                                                                                
assign out[5] = in[250];                                                                                                                                                                                                                                
assign out[6] = in[249];                                                                                                                                                                                                                                
assign out[7] = in[248];                                                                                                                                                                                                                                
assign out[8] = in[247];                                                                                                                                                                                                                                
assign out[9] = in[246];                                                                                                                                                                                                                                
assign out[10] = in[245];                                                                                                                                                                                                                               
assign out[11] = in[244];                                                                                                                                                                                                                               
assign out[12] = in[243];                                                                                                                                                                                                                               
assign out[13] = in[242];                                                                                                                                                                                                                               
assign out[14] = in[241];                                                                                                                                                                                                                               
assign out[15] = in[240];                                                                                                                                                                                                                               
assign out[16] = in[239];                                                                                                                                                                                                                               
assign out[17] = in[238];                                                                                                                                                                                                                               
assign out[18] = in[237];                                                                                                                                                                                                                               
assign out[19] = in[236];                                                                                                                                                                                                                               
assign out[20] = in[235];                                                                                                                                                                                                                               
assign out[21] = in[234];                                                                                                                                                                                                                               
assign out[22] = in[233];                                                                                                                                                                                                                               
assign out[23] = in[232];                                                                                                                                                                                                                               
assign out[24] = in[231];                                                                                                                                                                                                                               
assign out[25] = in[230];                                                                                                                                                                                                                               
assign out[26] = in[229];                                                                                                                                                                                                                               
assign out[27] = in[228];                                                                                                                                                                                                                               
assign out[28] = in[227];                                                                                                                                                                                                                               
assign out[29] = in[226];                                                                                                                                                                                                                               
assign out[30] = in[225];
assign out[31] = in[224];                                                                                                                                                                                                                               
assign out[32] = in[223];                                                                                                                                                                                                                               
assign out[33] = in[222];                                                                                                                                                                                                                               
assign out[34] = in[221];                                                                                                                                                                                                                               
assign out[35] = in[220];                                                                                                                                                                                                                               
assign out[36] = in[219];                                                                                                                                                                                                                               
assign out[37] = in[218];                                                                                                                                                                                                                               
assign out[38] = in[217];                                                                                                                                                                                                                               
assign out[39] = in[216];                                                                                                                                                                                                                               
assign out[40] = in[215];                                                                                                                                                                                                                               
assign out[41] = in[214];                                                                                                                                                                                                                               
assign out[42] = in[213];                                                                                                                                                                                                                               
assign out[43] = in[212];                                                                                                                                                                                                                               
assign out[44] = in[211];                                                                                                                                                                                                                               
assign out[45] = in[210];                                                                                                                                                                                                                               
assign out[46] = in[209];                                                                                                                                                                                                                               
assign out[47] = in[208];                                                                                                                                                                                                                               
assign out[48] = in[207];                                                                                                                                                                                                                               
assign out[49] = in[206];                                                                                                                                                                                                                               
assign out[50] = in[205];                                                                                                                                                                                                                               
assign out[51] = in[204];                                                                                                                                                                                                                               
assign out[52] = in[203];                                                                                                                                                                                                                               
assign out[53] = in[202];                                                                                                                                                                                                                               
assign out[54] = in[201];                                                                                                                                                                                                                               
assign out[55] = in[200];                                                                                                                                                                                                                               
assign out[56] = in[199];                                                                                                                                                                                                                               
assign out[57] = in[198];                                                                                                                                                                                                                               
assign out[58] = in[197];                                                                                                                                                                                                                               
assign out[59] = in[196];                                                                                                                                                                                                                               
assign out[60] = in[195];                                                                                                                                                                                                                               
assign out[61] = in[194];                                                                                                                                                                                                                               
assign out[62] = in[193];                                                                                                                                                                                                                               
assign out[63] = in[192];                                                                                                                                                                                                                               
assign out[64] = in[191];                                                                                                                                                                                                                               
assign out[65] = in[190];                                                                                                                                                                                                                               
assign out[66] = in[189];                                                                                                                                                                                                                               
assign out[67] = in[188];                                                                                                                                                                                                                               
assign out[68] = in[187];                                                                                                                                                                                                                               
assign out[69] = in[186];                                                                                                                                                                                                                               
assign out[70] = in[185];                                                                                                                                                                                                                               
assign out[71] = in[184];                                                                                                                                                                                                                               
assign out[72] = in[183];                                                                                                                                                                                                                               
assign out[73] = in[182];                                                                                                                                                                                                                               
assign out[74] = in[181];                                                                                                                                                                                                                               
assign out[75] = in[180];
assign out[76] = in[179];                                                                                                                                                                                                                               
assign out[77] = in[178];                                                                                                                                                                                                                               
assign out[78] = in[177];                                                                                                                                                                                                                               
assign out[79] = in[176];                                                                                                                                                                                                                               
assign out[80] = in[175];                                                                                                                                                                                                                               
assign out[81] = in[174];                                                                                                                                                                                                                               
assign out[82] = in[173];                                                                                                                                                                                                                               
assign out[83] = in[172];                                                                                                                                                                                                                               
assign out[84] = in[171];                                                                                                                                                                                                                               
assign out[85] = in[170];                                                                                                                                                                                                                               
assign out[86] = in[169];                                                                                                                                                                                                                               
assign out[87] = in[168];                                                                                                                                                                                                                               
assign out[88] = in[167];                                                                                                                                                                                                                               
assign out[89] = in[166];                                                                                                                                                                                                                               
assign out[90] = in[165];                                                                                                                                                                                                                               
assign out[91] = in[164];                                                                                                                                                                                                                               
assign out[92] = in[163];                                                                                                                                                                                                                               
assign out[93] = in[162];                                                                                                                                                                                                                               
assign out[94] = in[161];                                                                                                                                                                                                                               
assign out[95] = in[160];                                                                                                                                                                                                                               
assign out[96] = in[159];                                                                                                                                                                                                                               
assign out[97] = in[158];                                                                                                                                                                                                                               
assign out[98] = in[157];                                                                                                                                                                                                                               
assign out[99] = in[156];                                                                                                                                                                                                                               
assign out[100] = in[155];                                                                                                                                                                                                                              
assign out[101] = in[154];                                                                                                                                                                                                                              
assign out[102] = in[153];                                                                                                                                                                                                                              
assign out[103] = in[152];                                                                                                                                                                                                                              
assign out[104] = in[151];                                                                                                                                                                                                                              
assign out[105] = in[150];                                                                                                                                                                                                                              
assign out[106] = in[149];                                                                                                                                                                                                                              
assign out[107] = in[148];                                                                                                                                                                                                                              
assign out[108] = in[147];                                                                                                                                                                                                                              
assign out[109] = in[146];                                                                                                                                                                                                                              
assign out[110] = in[145];                                                                                                                                                                                                                              
assign out[111] = in[144];                                                                                                                                                                                                                              
assign out[112] = in[143];                                                                                                                                                                                                                              
assign out[113] = in[142];                                                                                                                                                                                                                              
assign out[114] = in[141];                                                                                                                                                                                                                              
assign out[115] = in[140];                                                                                                                                                                                                                              
assign out[116] = in[139];                                                                                                                                                                                                                              
assign out[117] = in[138];                                                                                                                                                                                                                              
assign out[118] = in[137];                                                                                                                                                                                                                              
assign out[119] = in[136];                                                                                                                                                                                                                              
assign out[120] = in[135];
assign out[121] = in[134];                                                                                                                                                                                                                              
assign out[122] = in[133];                                                                                                                                                                                                                              
assign out[123] = in[132];                                                                                                                                                                                                                              
assign out[124] = in[131];                                                                                                                                                                                                                              
assign out[125] = in[130];                                                                                                                                                                                                                              
assign out[126] = in[129];                                                                                                                                                                                                                              
assign out[127] = in[128];                                                                                                                                                                                                                              
assign out[128] = in[127];                                                                                                                                                                                                                              
assign out[129] = in[126];                                                                                                                                                                                                                              
assign out[130] = in[125];                                                                                                                                                                                                                              
assign out[131] = in[124];                                                                                                                                                                                                                              
assign out[132] = in[123];                                                                                                                                                                                                                              
assign out[133] = in[122];                                                                                                                                                                                                                              
assign out[134] = in[121];                                                                                                                                                                                                                              
assign out[135] = in[120];                                                                                                                                                                                                                              
assign out[136] = in[119];                                                                                                                                                                                                                              
assign out[137] = in[118];                                                                                                                                                                                                                              
assign out[138] = in[117];                                                                                                                                                                                                                              
assign out[139] = in[116];                                                                                                                                                                                                                              
assign out[140] = in[115];                                                                                                                                                                                                                              
assign out[141] = in[114];                                                                                                                                                                                                                              
assign out[142] = in[113];                                                                                                                                                                                                                              
assign out[143] = in[112];                                                                                                                                                                                                                              
assign out[144] = in[111];                                                                                                                                                                                                                              
assign out[145] = in[110];                                                                                                                                                                                                                              
assign out[146] = in[109];                                                                                                                                                                                                                              
assign out[147] = in[108];                                                                                                                                                                                                                              
assign out[148] = in[107];                                                                                                                                                                                                                              
assign out[149] = in[106];                                                                                                                                                                                                                              
assign out[150] = in[105];                                                                                                                                                                                                                              
assign out[151] = in[104];                                                                                                                                                                                                                              
assign out[152] = in[103];                                                                                                                                                                                                                              
assign out[153] = in[102];                                                                                                                                                                                                                              
assign out[154] = in[101];                                                                                                                                                                                                                              
assign out[155] = in[100];                                                                                                                                                                                                                              
assign out[156] = in[99];                                                                                                                                                                                                                               
assign out[157] = in[98];                                                                                                                                                                                                                               
assign out[158] = in[97];                                                                                                                                                                                                                               
assign out[159] = in[96];                                                                                                                                                                                                                               
assign out[160] = in[95];                                                                                                                                                                                                                               
assign out[161] = in[94];                                                                                                                                                                                                                               
assign out[162] = in[93];                                                                                                                                                                                                                               
assign out[163] = in[92];                                                                                                                                                                                                                               
assign out[164] = in[91];                                                                                                                                                                                                                               
assign out[165] = in[90];
assign out[166] = in[89];                                                                                                                                                                                                                               
assign out[167] = in[88];                                                                                                                                                                                                                               
assign out[168] = in[87];                                                                                                                                                                                                                               
assign out[169] = in[86];                                                                                                                                                                                                                               
assign out[170] = in[85];                                                                                                                                                                                                                               
assign out[171] = in[84];                                                                                                                                                                                                                               
assign out[172] = in[83];                                                                                                                                                                                                                               
assign out[173] = in[82];                                                                                                                                                                                                                               
assign out[174] = in[81];                                                                                                                                                                                                                               
assign out[175] = in[80];                                                                                                                                                                                                                               
assign out[176] = in[79];                                                                                                                                                                                                                               
assign out[177] = in[78];                                                                                                                                                                                                                               
assign out[178] = in[77];                                                                                                                                                                                                                               
assign out[179] = in[76];                                                                                                                                                                                                                               
assign out[180] = in[75];                                                                                                                                                                                                                               
assign out[181] = in[74];                                                                                                                                                                                                                               
assign out[182] = in[73];                                                                                                                                                                                                                               
assign out[183] = in[72];                                                                                                                                                                                                                               
assign out[184] = in[71];                                                                                                                                                                                                                               
assign out[185] = in[70];                                                                                                                                                                                                                               
assign out[186] = in[69];                                                                                                                                                                                                                               
assign out[187] = in[68];                                                                                                                                                                                                                               
assign out[188] = in[67];                                                                                                                                                                                                                               
assign out[189] = in[66];                                                                                                                                                                                                                               
assign out[190] = in[65];                                                                                                                                                                                                                               
assign out[191] = in[64];                                                                                                                                                                                                                               
assign out[192] = in[63];                                                                                                                                                                                                                               
assign out[193] = in[62];                                                                                                                                                                                                                               
assign out[194] = in[61];                                                                                                                                                                                                                               
assign out[195] = in[60];                                                                                                                                                                                                                               
assign out[196] = in[59];                                                                                                                                                                                                                               
assign out[197] = in[58];                                                                                                                                                                                                                               
assign out[198] = in[57];                                                                                                                                                                                                                               
assign out[199] = in[56];                                                                                                                                                                                                                               
assign out[200] = in[55];                                                                                                                                                                                                                               
assign out[201] = in[54];                                                                                                                                                                                                                               
assign out[202] = in[53];                                                                                                                                                                                                                               
assign out[203] = in[52];                                                                                                                                                                                                                               
assign out[204] = in[51];                                                                                                                                                                                                                               
assign out[205] = in[50];                                                                                                                                                                                                                               
assign out[206] = in[49];                                                                                                                                                                                                                               
assign out[207] = in[48];                                                                                                                                                                                                                               
assign out[208] = in[47];                                                                                                                                                                                                                               
assign out[209] = in[46];                                                                                                                                                                                                                               
assign out[210] = in[45];
assign out[211] = in[44];                                                                                                                                                                                                                               
assign out[212] = in[43];                                                                                                                                                                                                                               
assign out[213] = in[42];                                                                                                                                                                                                                               
assign out[214] = in[41];                                                                                                                                                                                                                               
assign out[215] = in[40];                                                                                                                                                                                                                               
assign out[216] = in[39];                                                                                                                                                                                                                               
assign out[217] = in[38];                                                                                                                                                                                                                               
assign out[218] = in[37];                                                                                                                                                                                                                               
assign out[219] = in[36];                                                                                                                                                                                                                               
assign out[220] = in[35];                                                                                                                                                                                                                               
assign out[221] = in[34];                                                                                                                                                                                                                               
assign out[222] = in[33];                                                                                                                                                                                                                               
assign out[223] = in[32];                                                                                                                                                                                                                               
assign out[224] = in[31];                                                                                                                                                                                                                               
assign out[225] = in[30];                                                                                                                                                                                                                               
assign out[226] = in[29];                                                                                                                                                                                                                               
assign out[227] = in[28];                                                                                                                                                                                                                               
assign out[228] = in[27];                                                                                                                                                                                                                               
assign out[229] = in[26];                                                                                                                                                                                                                               
assign out[230] = in[25];                                                                                                                                                                                                                               
assign out[231] = in[24];                                                                                                                                                                                                                               
assign out[232] = in[23];                                                                                                                                                                                                                               
assign out[233] = in[22];                                                                                                                                                                                                                               
assign out[234] = in[21];                                                                                                                                                                                                                               
assign out[235] = in[20];                                                                                                                                                                                                                               
assign out[236] = in[19];                                                                                                                                                                                                                               
assign out[237] = in[18];                                                                                                                                                                                                                               
assign out[238] = in[17];                                                                                                                                                                                                                               
assign out[239] = in[16];                                                                                                                                                                                                                               
assign out[240] = in[15];                                                                                                                                                                                                                               
assign out[241] = in[14];                                                                                                                                                                                                                               
assign out[242] = in[13];                                                                                                                                                                                                                               
assign out[243] = in[12];                                                                                                                                                                                                                               
assign out[244] = in[11];                                                                                                                                                                                                                               
assign out[245] = in[10];                                                                                                                                                                                                                               
assign out[246] = in[9];                                                                                                                                                                                                                                
assign out[247] = in[8];                                                                                                                                                                                                                                
assign out[248] = in[7];                                                                                                                                                                                                                                
assign out[249] = in[6];                                                                                                                                                                                                                                
assign out[250] = in[5];                                                                                                                                                                                                                                
assign out[251] = in[4];                                                                                                                                                                                                                                
assign out[252] = in[3];                                                                                                                                                                                                                                
assign out[253] = in[2];                                                                                                                                                                                                                                
assign out[254] = in[1];                                                                                                                                                                                                                                
assign out[255] = in[0];
endmodule
