module SHA256(in,out);
input [511:0]in;
output [255:0]out;
//64 k constants
parameter k1= 32'h428A2F98;
parameter k2 = 32'h71374491;
parameter k3 = 32'hB5C0FBCF;
parameter k4 = 32'hE9B5DBA5;
parameter k5 = 32'h3956C25B;
parameter k6 = 32'h59F111F1;
parameter k7 = 32'h923F82A4;
parameter k8 = 32'hAB1C5ED5;
parameter k9 = 32'hD807AA98;
parameter k10 = 32'h12835B01;
parameter k11 = 32'h243185BE;
parameter k12 = 32'h550C7DC3;
parameter k13 = 32'h72BE5D74;
parameter k14 = 32'h80DEB1FE;
parameter k15 = 32'h9BDC06A7;
parameter k16 = 32'hC19BF174;
parameter k17 = 32'hE49B69C1;
parameter k18 = 32'hEFBE4786;
parameter k19 = 32'h0FC19DC6;
parameter k20 = 32'h240CA1CC;
parameter k21 = 32'h2DE92C6F;
parameter k22 = 32'h4A7484AA;
parameter k23 = 32'h5CB0A9DC;
parameter k24 = 32'h76F988DA;
parameter k25 = 32'h983E5152;
parameter k26 = 32'hA831C66D;
parameter k27 = 32'hB00327C8;
parameter k28 = 32'hBF597FC7;
parameter k29 = 32'hC6E00BF3;
parameter k30 = 32'hD5A79147;
parameter k31 = 32'h06CA6351;
parameter k32 = 32'h14292967;
parameter k33 = 32'h27B70A85;
parameter k34 = 32'h2E1B2138;
parameter k35 = 32'h4D2C6DFC;
parameter k36 = 32'h53380D13;
parameter k37 = 32'h650A7354;
parameter k38 = 32'h766A0ABB;
parameter k39 = 32'h81C2C92E;
parameter k40 = 32'h92722C85;
parameter k41 = 32'hA2BFE8A1;
parameter k42 = 32'hA81A664B;
parameter k43 = 32'hC24B8B70;
parameter k44 = 32'hC76C51A3;
parameter k45 = 32'hD192E819;
parameter k46 = 32'hD6990624;
parameter k47 = 32'hF40E3585;
parameter k48 = 32'h106AA070;
parameter k49 = 32'h19A4C116;
parameter k50 = 32'h1E376C08;
parameter k51 = 32'h2748774C;
parameter k52 = 32'h34B0BCB5;
parameter k53 = 32'h391C0CB3;
parameter k54 = 32'h4ED8AA4A;
parameter k55 = 32'h5B9CCA4F;
parameter k56 = 32'h682E6FF3;
parameter k57 = 32'h748F82EE;
parameter k58 = 32'h78A5636F;
parameter k59 = 32'h84C87814;
parameter k60 = 32'h8CC70208;
parameter k61 = 32'h90BEFFFA;
parameter k62 = 32'hA4506CEB;
parameter k63 = 32'hBEF9A3F7;
parameter k64 = 32'hC67178F2;
wire [31:0]w1;
wire [31:0]w2;
wire [31:0]w3;
wire [31:0]w4;
wire [31:0]w5;
wire [31:0]w6;
wire [31:0]w7;
wire [31:0]w8;
wire [31:0]w9;
wire [31:0]w10;
wire [31:0]w11;
wire [31:0]w12;
wire [31:0]w13;
wire [31:0]w14;
wire [31:0]w15;
wire [31:0]w16;
wire [31:0]w17;
wire [31:0]w18;
wire [31:0]w19;
wire [31:0]w20;
wire [31:0]w21;
wire [31:0]w22;
wire [31:0]w23;
wire [31:0]w24;
wire [31:0]w25;
wire [31:0]w26;
wire [31:0]w27;
wire [31:0]w28;
wire [31:0]w29;
wire [31:0]w30;
wire [31:0]w31;
wire [31:0]w32;
wire [31:0]w33;
wire [31:0]w34;
wire [31:0]w35;
wire [31:0]w36;
wire [31:0]w37;
wire [31:0]w38;
wire [31:0]w39;
wire [31:0]w40;
wire [31:0]w41;
wire [31:0]w42;
wire [31:0]w43;
wire [31:0]w44;
wire [31:0]w45;
wire [31:0]w46;
wire [31:0]w47;
wire [31:0]w48;
wire [31:0]w49;
wire [31:0]w50;
wire [31:0]w51;
wire [31:0]w52;
wire [31:0]w53;
wire [31:0]w54;
wire [31:0]w55;
wire [31:0]w56;
wire [31:0]w57;
wire [31:0]w58;
wire [31:0]w59;
wire [31:0]w60;
wire [31:0]w61;
wire [31:0]w62;
wire [31:0]w63;
wire [31:0]w64;
wire [31:0]aout;
wire [31:0]bout;
wire [31:0]cout;
wire [31:0]dout;
wire [31:0]eout;
wire [31:0]fout;
wire [31:0]gout;
wire [31:0]hout;
//initial constants
parameter ainit= 32'h6A09E667;
parameter binit= 32'hBB67AE85;
parameter cinit= 32'h3C6EF372;
parameter dinit= 32'hA54FF53A;
parameter einit= 32'h510E527F;
parameter finit= 32'h9B05688C;
parameter ginit= 32'h1F83D9AB;
parameter hinit= 32'h5BE0CD19;
//prenodes w assignments
assign w1=in[511:480];
assign w2=in[479:448];
assign w3=in[447:416];
assign w4=in[414:384];
assign w5=in[383:352];
assign w6=in[351:320];
assign w7=in[319:288];
assign w8=in[287:256];
assign w9=in[255:224];
assign w10=in[223:192];
assign w11=in[191:160];
assign w12=in[159:128];
assign w13=in[127:96];
assign w14=in[95:64];
assign w15=in[63:32];
assign w16=in[31:0];
wassign was17(w2,w15,w1,w10,w17);
wassign was18(w3,w16,w2,w11,w18);
wassign was19(w4,w17,w3,w12,w19);
wassign was20(w5,w18,w4,w13,w20);
wassign was21(w6,w19,w5,w14,w21);
wassign was22(w7,w20,w6,w15,w22);
wassign was23(w8,w21,w7,w16,w23);
wassign was24(w9,w22,w8,w17,w24);
wassign was25(w10,w23,w9,w18,w25);
wassign was26(w11,w24,w10,w19,w26);
wassign was27(w12,w25,w11,w20,w27);
wassign was28(w13,w26,w12,w21,w28);
wassign was29(w14,w27,w13,w22,w29);
wassign was30(w15,w28,w14,w23,w30);
wassign was31(w16,w29,w15,w24,w31);
wassign was32(w17,w30,w16,w25,w32);
wassign was33(w18,w31,w17,w26,w33);
wassign was34(w19,w32,w18,w27,w34);
wassign was35(w20,w33,w19,w28,w35);
wassign was36(w21,w34,w20,w29,w36);
wassign was37(w22,w35,w21,w30,w37);
wassign was38(w23,w36,w22,w31,w38);
wassign was39(w24,w37,w23,w32,w39);
wassign was40(w25,w38,w24,w33,w40);
wassign was41(w26,w39,w25,w34,w41);
wassign was42(w27,w40,w26,w35,w42);
wassign was43(w28,w41,w27,w36,w43);
wassign was44(w29,w42,w28,w37,w44);
wassign was45(w30,w43,w29,w38,w45);
wassign was46(w31,w44,w30,w39,w46);
wassign was47(w32,w45,w31,w40,w47);
wassign was48(w33,w46,w32,w41,w48);
wassign was49(w34,w47,w33,w42,w49);
wassign was50(w35,w48,w34,w43,w50);
wassign was51(w36,w49,w35,w44,w51);
wassign was52(w37,w50,w36,w45,w52);
wassign was53(w38,w51,w37,w46,w53);
wassign was54(w39,w52,w38,w47,w54);
wassign was55(w40,w53,w39,w48,w55);
wassign was56(w41,w54,w40,w49,w56);
wassign was57(w42,w55,w41,w50,w57);
wassign was58(w43,w56,w42,w51,w58);
wassign was59(w44,w57,w43,w52,w59);
wassign was60(w45,w58,w44,w53,w60);
wassign was61(w46,w59,w45,w54,w61);
wassign was62(w47,w60,w46,w55,w62);
wassign was63(w48,w61,w47,w56,w63);
wassign was64(w49,w62,w48,w57,w64);
//begins 64 cycles of hashing
wire [31:0]a1;
wire [31:0]b1;
wire [31:0]c1;
wire [31:0]d1;
wire [31:0]e1;
wire [31:0]f1;
wire [31:0]g1;
wire [31:0]h1;
SHA256Node node1(ainit,binit,cinit,dinit,einit,finit,ginit,hinit,a1,b1,c1,d1,e1,f1,g1,h1,k1,w1);
wire [31:0]a2;                                                                                                                                                                                                                                         
wire [31:0]b2;                                                                                                                                                                                                                                         
wire [31:0]c2;                                                                                                                                                                                                                                         
wire [31:0]d2;                                                                                                                                                                                                                                         
wire [31:0]e2;                                                                                                                                                                                                                                         
wire [31:0]f2;                                                                                                                                                                                                                                         
wire [31:0]g2;
wire [31:0]h2;                                                                                                                                                                                                                                         
SHA256Node node2(a1,b1,c1,d1,e1,f1,g1,h1,a2,b2,c2,d2,e2,f2,g2,h2,k2,w2);
wire [31:0]a3;                                                                                                                                                                                                                                         
wire [31:0]b3;                                                                                                                                                                                                                                         
wire [31:0]c3;                                                                                                                                                                                                                                         
wire [31:0]d3;                                                                                                                                                                                                                                         
wire [31:0]e3;                                                                                                                                                                                                                                         
wire [31:0]f3;                                                                                                                                                                                                                                         
wire [31:0]g3;
wire [31:0]h3;                                                                                                                                                                                                                                         
SHA256Node node3(a2,b2,c2,d2,e2,f2,g2,h2,a3,b3,c3,d3,e3,f3,g3,h3,k3,w3);
wire [31:0]a4;                                                                                                                                                                                                                                         
wire [31:0]b4;                                                                                                                                                                                                                                         
wire [31:0]c4;                                                                                                                                                                                                                                         
wire [31:0]d4;                                                                                                                                                                                                                                         
wire [31:0]e4;                                                                                                                                                                                                                                         
wire [31:0]f4;                                                                                                                                                                                                                                         
wire [31:0]g4;
wire [31:0]h4;                                                                                                                                                                                                                                         
SHA256Node node4(a3,b3,c3,d3,e3,f3,g3,h3,a4,b4,c4,d4,e4,f4,g4,h4,k4,w4);
wire [31:0]a5;                                                                                                                                                                                                                                         
wire [31:0]b5;                                                                                                                                                                                                                                         
wire [31:0]c5;                                                                                                                                                                                                                                         
wire [31:0]d5;                                                                                                                                                                                                                                         
wire [31:0]e5;                                                                                                                                                                                                                                         
wire [31:0]f5;                                                                                                                                                                                                                                         
wire [31:0]g5;
wire [31:0]h5;                                                                                                                                                                                                                                         
SHA256Node node5(a4,b4,c4,d4,e4,f4,g4,h4,a5,b5,c5,d5,e5,f5,g5,h5,k5,w5);
wire [31:0]a6;                                                                                                                                                                                                                                          
wire [31:0]b6;                                                                                                                                                                                                                                          
wire [31:0]c6;                                                                                                                                                                                                                                          
wire [31:0]d6;                                                                                                                                                                                                                                          
wire [31:0]e6;                                                                                                                                                                                                                                          
wire [31:0]f6;                                                                                                                                                                                                                                          
wire [31:0]g6;
wire [31:0]h6;                                                                                                                                                                                                                                          
SHA256Node node6(a5,b5,c5,d5,e5,f5,g5,h5,a6,b6,c6,d6,e6,f6,g6,h6,k6,w6);                                                                                                                                                                                      
wire [31:0]a7;                                                                                                                                                                                                                                          
wire [31:0]b7;                                                                                                                                                                                                                                          
wire [31:0]c7;                                                                                                                                                                                                                                          
wire [31:0]d7;                                                                                                                                                                                                                                          
wire [31:0]e7;                                                                                                                                                                                                                                          
wire [31:0]f7;                                                                                                                                                                                                                                          
wire [31:0]g7;
wire [31:0]h7;                                                                                                                                                                                                                                          
SHA256Node node7(a6,b6,c6,d6,e6,f6,g6,h6,a7,b7,c7,d7,e7,f7,g7,h7,k7,w7);                                                                                                                                                                                      
wire [31:0]a8;                                                                                                                                                                                                                                          
wire [31:0]b8;                                                                                                                                                                                                                                          
wire [31:0]c8;                                                                                                                                                                                                                                          
wire [31:0]d8;                                                                                                                                                                                                                                          
wire [31:0]e8;                                                                                                                                                                                                                                          
wire [31:0]f8;                                                                                                                                                                                                                                          
wire [31:0]g8;
wire [31:0]h8;                                                                                                                                                                                                                                          
SHA256Node node8(a7,b7,c7,d7,e7,f7,g7,h7,a8,b8,c8,d8,e8,f8,g8,h8,k8,w8);                                                                                                                                                                                      
wire [31:0]a9;                                                                                                                                                                                                                                          
wire [31:0]b9;                                                                                                                                                                                                                                          
wire [31:0]c9;                                                                                                                                                                                                                                          
wire [31:0]d9;                                                                                                                                                                                                                                          
wire [31:0]e9;                                                                                                                                                                                                                                          
wire [31:0]f9;                                                                                                                                                                                                                                          
wire [31:0]g9;
wire [31:0]h9;                                                                                                                                                                                                                                          
SHA256Node node9(a8,b8,c8,d8,e8,f8,g8,h8,a9,b9,c9,d9,e9,f9,g9,h9,k9,w9);
wire [31:0]a10;                                                                                                                                                                                                                                         
wire [31:0]b10;                                                                                                                                                                                                                                         
wire [31:0]c10;                                                                                                                                                                                                                                         
wire [31:0]d10;                                                                                                                                                                                                                                         
wire [31:0]e10;                                                                                                                                                                                                                                         
wire [31:0]f10;                                                                                                                                                                                                                                         
wire [31:0]g10;
wire [31:0]h10;                                                                                                                                                                                                                                         
SHA256Node node10(a9,b9,c9,d9,e9,f9,g9,h10,a10,b10,c10,d10,e10,f10,g10,h10,k10,w10);                                                                                                                                                                            
wire [31:0]a11;                                                                                                                                                                                                                                         
wire [31:0]b11;                                                                                                                                                                                                                                         
wire [31:0]c11;                                                                                                                                                                                                                                         
wire [31:0]d11;                                                                                                                                                                                                                                         
wire [31:0]e11;                                                                                                                                                                                                                                         
wire [31:0]f11;                                                                                                                                                                                                                                         
wire [31:0]g11;
wire [31:0]h11;                                                                                                                                                                                                                                         
SHA256Node node11(a10,b10,c10,d10,e10,f10,g10,h10,a11,b11,c11,d11,e11,f11,g11,h11,k11,w11);                                                                                                                                                                     
wire [31:0]a12;                                                                                                                                                                                                                                         
wire [31:0]b12;                                                                                                                                                                                                                                         
wire [31:0]c12;                                                                                                                                                                                                                                         
wire [31:0]d12;                                                                                                                                                                                                                                         
wire [31:0]e12;                                                                                                                                                                                                                                         
wire [31:0]f12;                                                                                                                                                                                                                                         
wire [31:0]g12;
wire [31:0]h12;                                                                                                                                                                                                                                         
SHA256Node node12(a11,b11,c11,d11,e11,f11,g11,h11,a12,b12,c12,d12,e12,f12,g12,h12,k12,w12);                                                                                                                                                                     
wire [31:0]a13;                                                                                                                                                                                                                                         
wire [31:0]b13;                                                                                                                                                                                                                                         
wire [31:0]c13;                                                                                                                                                                                                                                         
wire [31:0]d13;                                                                                                                                                                                                                                         
wire [31:0]e13;                                                                                                                                                                                                                                         
wire [31:0]f13;                                                                                                                                                                                                                                         
wire [31:0]g13;
wire [31:0]h13;                                                                                                                                                                                                                                         
SHA256Node node13(a12,b12,c12,d12,e12,f12,g12,h12,a13,b13,c13,d13,e13,f13,g13,h13,k13,w13);                                                                                                                                                                     
wire [31:0]a14;                                                                                                                                                                                                                                         
wire [31:0]b14;                                                                                                                                                                                                                                         
wire [31:0]c14;                                                                                                                                                                                                                                         
wire [31:0]d14;                                                                                                                                                                                                                                         
wire [31:0]e14;                                                                                                                                                                                                                                         
wire [31:0]f14;                                                                                                                                                                                                                                         
wire [31:0]g14;
wire [31:0]h14;                                                                                                                                                                                                                                         
SHA256Node node14(a13,b13,c13,d13,e13,f13,g13,h13,a14,b14,c14,d14,e14,f14,g14,h14,k14,w14);
wire [31:0]a15;                                                                                                                                                                                                                                         
wire [31:0]b15;                                                                                                                                                                                                                                         
wire [31:0]c15;                                                                                                                                                                                                                                         
wire [31:0]d15;                                                                                                                                                                                                                                         
wire [31:0]e15;                                                                                                                                                                                                                                         
wire [31:0]f15;                                                                                                                                                                                                                                         
wire [31:0]g15;
wire [31:0]h15;                                                                                                                                                                                                                                         
SHA256Node node15(a14,b14,c14,d14,e14,f14,g14,h14,a15,b15,c15,d15,e15,f15,g15,h15,k15,w15);                                                                                                                                                                     
wire [31:0]a16;                                                                                                                                                                                                                                         
wire [31:0]b16;                                                                                                                                                                                                                                         
wire [31:0]c16;                                                                                                                                                                                                                                         
wire [31:0]d16;                                                                                                                                                                                                                                         
wire [31:0]e16;                                                                                                                                                                                                                                         
wire [31:0]f16;                                                                                                                                                                                                                                         
wire [31:0]g16;
wire [31:0]h16;                                                                                                                                                                                                                                         
SHA256Node node16(a15,b15,c15,d15,e15,f15,g15,h15,a16,b16,c16,d16,e16,f16,g16,h16,k16,w16);                                                                                                                                                                     
wire [31:0]a17;                                                                                                                                                                                                                                         
wire [31:0]b17;                                                                                                                                                                                                                                         
wire [31:0]c17;                                                                                                                                                                                                                                         
wire [31:0]d17;                                                                                                                                                                                                                                         
wire [31:0]e17;                                                                                                                                                                                                                                         
wire [31:0]f17;                                                                                                                                                                                                                                         
wire [31:0]g17;
wire [31:0]h17;                                                                                                                                                                                                                                         
SHA256Node node17(a16,b16,c16,d16,e16,f16,g16,h16,a17,b17,c17,d17,e17,f17,g17,h17,k17,w17);                                                                                                                                                                     
wire [31:0]a18;                                                                                                                                                                                                                                         
wire [31:0]b18;                                                                                                                                                                                                                                         
wire [31:0]c18;                                                                                                                                                                                                                                         
wire [31:0]d18;                                                                                                                                                                                                                                         
wire [31:0]e18;                                                                                                                                                                                                                                         
wire [31:0]f18;                                                                                                                                                                                                                                         
wire [31:0]g18;
wire [31:0]h18;                                                                                                                                                                                                                                         
SHA256Node node18(a17,b17,c17,d17,e17,f17,g17,h17,a18,b18,c18,d18,e18,f18,g18,h18,k18,w18);                                                                                                                                                                     
wire [31:0]a19;                                                                                                                                                                                                                                         
wire [31:0]b19;                                                                                                                                                                                                                                         
wire [31:0]c19;                                                                                                                                                                                                                                         
wire [31:0]d19;                                                                                                                                                                                                                                         
wire [31:0]e19;                                                                                                                                                                                                                                         
wire [31:0]f19;                                                                                                                                                                                                                                         
wire [31:0]g19;
wire [31:0]h19;                                                                                                                                                                                                                                         
SHA256Node node19(a18,b18,c18,d18,e18,f18,g18,h18,a19,b19,c19,d19,e19,f19,g19,h19,k19,w19);
wire [31:0]a20;                                                                                                                                                                                                                                         
wire [31:0]b20;                                                                                                                                                                                                                                         
wire [31:0]c20;                                                                                                                                                                                                                                         
wire [31:0]d20;                                                                                                                                                                                                                                         
wire [31:0]e20;                                                                                                                                                                                                                                         
wire [31:0]f20;                                                                                                                                                                                                                                         
wire [31:0]g20;
wire [31:0]h20;                                                                                                                                                                                                                                         
SHA256Node node20(a19,b19,c19,d19,e19,f19,g19,h19,a20,b20,c20,d20,e20,f20,g20,h20,k20,w20);                                                                                                                                                                     
wire [31:0]a21;                                                                                                                                                                                                                                         
wire [31:0]b21;                                                                                                                                                                                                                                         
wire [31:0]c21;                                                                                                                                                                                                                                         
wire [31:0]d21;                                                                                                                                                                                                                                         
wire [31:0]e21;                                                                                                                                                                                                                                         
wire [31:0]f21;                                                                                                                                                                                                                                         
wire [31:0]g21;
wire [31:0]h21;                                                                                                                                                                                                                                         
SHA256Node node21(a20,b20,c20,d20,e20,f20,g20,h20,a21,b21,c21,d21,e21,f21,g21,h21,k21,w21);                                                                                                                                                                     
wire [31:0]a22;                                                                                                                                                                                                                                         
wire [31:0]b22;                                                                                                                                                                                                                                         
wire [31:0]c22;                                                                                                                                                                                                                                         
wire [31:0]d22;                                                                                                                                                                                                                                         
wire [31:0]e22;                                                                                                                                                                                                                                         
wire [31:0]f22;                                                                                                                                                                                                                                         
wire [31:0]g22;
wire [31:0]h22;                                                                                                                                                                                                                                         
SHA256Node node22(a21,b21,c21,d21,e21,f21,g21,h21,a22,b22,c22,d22,e22,f22,g22,h22,k22,w22);                                                                                                                                                                     
wire [31:0]a23;                                                                                                                                                                                                                                         
wire [31:0]b23;                                                                                                                                                                                                                                         
wire [31:0]c23;                                                                                                                                                                                                                                         
wire [31:0]d23;                                                                                                                                                                                                                                         
wire [31:0]e23;                                                                                                                                                                                                                                         
wire [31:0]f23;                                                                                                                                                                                                                                         
wire [31:0]g23;
wire [31:0]h23;                                                                                                                                                                                                                                        
SHA256Node node23(a22,b22,c22,d22,e22,f22,g22,h22,a23,b23,c23,d23,e23,f23,g23,h23,k23,w23);                                                                                                                                                                     
wire [31:0]a24;                                                                                                                                                                                                                                         
wire [31:0]b24;                                                                                                                                                                                                                                         
wire [31:0]c24;                                                                                                                                                                                                                                         
wire [31:0]d24;                                                                                                                                                                                                                                         
wire [31:0]e24;                                                                                                                                                                                                                                         
wire [31:0]f24;                                                                                                                                                                                                                                         
wire [31:0]g24;
wire [31:0]h24;                                                                                                                                                                                                                                         
SHA256Node node24(a23,b23,c23,d23,e23,f23,g23,h23,a24,b24,c24,d24,e24,f24,g24,h24,k24,w24);
wire [31:0]a25;                                                                                                                                                                                                                                         
wire [31:0]b25;                                                                                                                                                                                                                                         
wire [31:0]c25;                                                                                                                                                                                                                                         
wire [31:0]d25;                                                                                                                                                                                                                                         
wire [31:0]e25;                                                                                                                                                                                                                                         
wire [31:0]f25;                                                                                                                                                                                                                                         
wire [31:0]g25;
wire [31:0]h25;                                                                                                                                                                                                                                         
SHA256Node node25(a24,b24,c24,d24,e24,f24,g24,h24,a25,b25,c25,d25,e25,f25,g25,h25,k25,w25);                                                                                                                                                                     
wire [31:0]a26;                                                                                                                                                                                                                                         
wire [31:0]b26;                                                                                                                                                                                                                                         
wire [31:0]c26;                                                                                                                                                                                                                                         
wire [31:0]d26;                                                                                                                                                                                                                                         
wire [31:0]e26;                                                                                                                                                                                                                                         
wire [31:0]f26;                                                                                                                                                                                                                                         
wire [31:0]g26;
wire [31:0]h26;                                                                                                                                                                                                                                         
SHA256Node node26(a25,b25,c25,d25,e25,f25,g25,h25,a26,b26,c26,d26,e26,f26,g26,h26,k26,w26);                                                                                                                                                                     
wire [31:0]a27;                                                                                                                                                                                                                                         
wire [31:0]b27;                                                                                                                                                                                                                                         
wire [31:0]c27;                                                                                                                                                                                                                                         
wire [31:0]d27;                                                                                                                                                                                                                                         
wire [31:0]e27;                                                                                                                                                                                                                                         
wire [31:0]f27;                                                                                                                                                                                                                                         
wire [31:0]g27;
wire [31:0]h27;                                                                                                                                                                                                                                         
SHA256Node node27(a26,b26,c26,d26,e26,f26,g26,h26,a27,b27,c27,d27,e27,f27,g27,h27,k27,w27);                                                                                                                                                                     
wire [31:0]a28;                                                                                                                                                                                                                                         
wire [31:0]b28;                                                                                                                                                                                                                                         
wire [31:0]c28;                                                                                                                                                                                                                                         
wire [31:0]d28;                                                                                                                                                                                                                                         
wire [31:0]e28;                                                                                                                                                                                                                                         
wire [31:0]f28;                                                                                                                                                                                                                                         
wire [31:0]g28;
wire [31:0]h28;                                                                                                                                                                                                                                         
SHA256Node node28(a27,b27,c27,d27,e27,f27,g27,h27,a28,b28,c28,d28,e28,f28,g28,h28,k28,w28);                                                                                                                                                                     
wire [31:0]a29;                                                                                                                                                                                                                                         
wire [31:0]b29;                                                                                                                                                                                                                                         
wire [31:0]c29;                                                                                                                                                                                                                                         
wire [31:0]d29;                                                                                                                                                                                                                                         
wire [31:0]e29;                                                                                                                                                                                                                                         
wire [31:0]f29;                                                                                                                                                                                                                                         
wire [31:0]g29;
wire [31:0]h29;                                                                                                                                                                                                                                         
SHA256Node node29(a28,b28,c28,d28,e28,f28,g28,h28,a29,b29,c29,d29,e29,f29,g29,h29,k29,w29);
wire [31:0]a30;                                                                                                                                                                                                                                         
wire [31:0]b30;                                                                                                                                                                                                                                         
wire [31:0]c30;                                                                                                                                                                                                                                         
wire [31:0]d30;                                                                                                                                                                                                                                         
wire [31:0]e30;                                                                                                                                                                                                                                         
wire [31:0]f30;                                                                                                                                                                                                                                         
wire [31:0]g30;
wire [31:0]h30;                                                                                                                                                                                                                                         
SHA256Node node30(a29,b29,c29,d29,e29,f29,g29,h29,a30,b30,c30,d30,e30,f30,g30,h30,k30,w30);                                                                                                                                                                     
wire [31:0]a31;                                                                                                                                                                                                                                         
wire [31:0]b31;                                                                                                                                                                                                                                         
wire [31:0]c31;                                                                                                                                                                                                                                         
wire [31:0]d31;                                                                                                                                                                                                                                         
wire [31:0]e31;                                                                                                                                                                                                                                         
wire [31:0]f31;                                                                                                                                                                                                                                         
wire [31:0]g31;
wire [31:0]h31;                                                                                                                                                                                                                                         
SHA256Node node31(a30,b30,c30,d30,e30,f30,g30,h30,a31,b31,c31,d31,e31,f31,g31,h31,k31,w31);                                                                                                                                                                     
wire [31:0]a32;                                                                                                                                                                                                                                         
wire [31:0]b32;                                                                                                                                                                                                                                         
wire [31:0]c32;                                                                                                                                                                                                                                         
wire [31:0]d32;                                                                                                                                                                                                                                         
wire [31:0]e32;                                                                                                                                                                                                                                         
wire [31:0]f32;                                                                                                                                                                                                                                         
wire [31:0]g32;
wire [31:0]h32;                                                                                                                                                                                                                                         
SHA256Node node32(a31,b31,c31,d31,e31,f31,g31,h31,a32,b32,c32,d32,e32,f32,g32,h32,k32,w32);                                                                                                                                                                     
wire [31:0]a33;                                                                                                                                                                                                                                         
wire [31:0]b33;                                                                                                                                                                                                                                         
wire [31:0]c33;                                                                                                                                                                                                                                         
wire [31:0]d33;                                                                                                                                                                                                                                         
wire [31:0]e33;                                                                                                                                                                                                                                         
wire [31:0]f33;                                                                                                                                                                                                                                         
wire [31:0]g33;
wire [31:0]h33;                                                                                                                                                                                                                                         
SHA256Node node33(a32,b32,c32,d32,e32,f32,g32,h32,a33,b33,c33,d33,e33,f33,g33,h33,k33,w33);                                                                                                                                                                     
wire [31:0]a34;                                                                                                                                                                                                                                         
wire [31:0]b34;                                                                                                                                                                                                                                         
wire [31:0]c34;                                                                                                                                                                                                                                         
wire [31:0]d34;                                                                                                                                                                                                                                         
wire [31:0]e34;                                                                                                                                                                                                                                         
wire [31:0]f34;                                                                                                                                                                                                                                         
wire [31:0]g34;
wire [31:0]h34;                                                                                                                                                                                                                                         
SHA256Node node34(a33,b33,c33,d33,e33,f33,g33,h33,a34,b34,c34,d34,e34,f34,g34,h34,k34,w34);
wire [31:0]a35;                                                                                                                                                                                                                                         
wire [31:0]b35;                                                                                                                                                                                                                                         
wire [31:0]c35;                                                                                                                                                                                                                                         
wire [31:0]d35;                                                                                                                                                                                                                                         
wire [31:0]e35;                                                                                                                                                                                                                                         
wire [31:0]f35;                                                                                                                                                                                                                                         
wire [31:0]g35;
wire [31:0]h35;                                                                                                                                                                                                                                         
SHA256Node node35(a34,b34,c34,d34,e34,f34,g34,h34,a35,b35,c35,d35,e35,f35,g35,h35,k35,w35);                                                                                                                                                                     
wire [31:0]a36;                                                                                                                                                                                                                                         
wire [31:0]b36;                                                                                                                                                                                                                                         
wire [31:0]c36;                                                                                                                                                                                                                                         
wire [31:0]d36;                                                                                                                                                                                                                                         
wire [31:0]e36;                                                                                                                                                                                                                                         
wire [31:0]f36;                                                                                                                                                                                                                                         
wire [31:0]g36;
wire [31:0]h36;                                                                                                                                                                                                                                         
SHA256Node node36(a35,b35,c35,d35,e35,f35,g35,h35,a36,b36,c36,d36,e36,f36,g36,h36,k36,w36);                                                                                                                                                                     
wire [31:0]a37;                                                                                                                                                                                                                                         
wire [31:0]b37;                                                                                                                                                                                                                                         
wire [31:0]c37;                                                                                                                                                                                                                                         
wire [31:0]d37;                                                                                                                                                                                                                                         
wire [31:0]e37;                                                                                                                                                                                                                                         
wire [31:0]f37;                                                                                                                                                                                                                                         
wire [31:0]g37;
wire [31:0]h37;                                                                                                                                                                                                                                         
SHA256Node node37(a36,b36,c36,d36,e36,f36,g36,h36,a37,b37,c37,d37,e37,f37,g37,h37,k37,w37);                                                                                                                                                                     
wire [31:0]a38;                                                                                                                                                                                                                                         
wire [31:0]b38;                                                                                                                                                                                                                                         
wire [31:0]c38;                                                                                                                                                                                                                                         
wire [31:0]d38;                                                                                                                                                                                                                                         
wire [31:0]e38;                                                                                                                                                                                                                                         
wire [31:0]f38;                                                                                                                                                                                                                                         
wire [31:0]g38;
wire [31:0]h38;                                                                                                                                                                                                                                         
SHA256Node node38(a37,b37,c37,d37,e37,f37,g37,h37,a38,b38,c38,d38,e38,f38,g38,h38,k38,w38);                                                                                                                                                                     
wire [31:0]a39;                                                                                                                                                                                                                                         
wire [31:0]b39;                                                                                                                                                                                                                                         
wire [31:0]c39;                                                                                                                                                                                                                                         
wire [31:0]d39;                                                                                                                                                                                                                                         
wire [31:0]e39;                                                                                                                                                                                                                                         
wire [31:0]f39;                                                                                                                                                                                                                                         
wire [31:0]g39;
wire [31:0]h39;                                                                                                                                                                                                                                         
SHA256Node node39(a38,b38,c38,d38,e38,f38,g38,h38,a39,b39,c39,d39,e39,f39,g39,h39,k39,w39);
wire [31:0]a40;                                                                                                                                                                                                                                         
wire [31:0]b40;                                                                                                                                                                                                                                         
wire [31:0]c40;                                                                                                                                                                                                                                         
wire [31:0]d40;                                                                                                                                                                                                                                         
wire [31:0]e40;                                                                                                                                                                                                                                         
wire [31:0]f40;                                                                                                                                                                                                                                         
wire [31:0]g40;
wire [31:0]h40;                                                                                                                                                                                                                                         
SHA256Node node40(a39,b39,c39,d39,e39,f39,g39,h39,a40,b40,c40,d40,e40,f40,g40,h40,k40,w40);                                                                                                                                                                     
wire [31:0]a41;                                                                                                                                                                                                                                         
wire [31:0]b41;                                                                                                                                                                                                                                         
wire [31:0]c41;                                                                                                                                                                                                                                         
wire [31:0]d41;                                                                                                                                                                                                                                         
wire [31:0]e41;                                                                                                                                                                                                                                         
wire [31:0]f41;                                                                                                                                                                                                                                         
wire [31:0]g41;
wire [31:0]h41;                                                                                                                                                                                                                                         
SHA256Node node41(a40,b40,c40,d40,e40,f40,g40,h40,a41,b41,c41,d41,e41,f41,g41,h41,k41,w41);                                                                                                                                                                     
wire [31:0]a42;                                                                                                                                                                                                                                         
wire [31:0]b42;                                                                                                                                                                                                                                         
wire [31:0]c42;                                                                                                                                                                                                                                         
wire [31:0]d42;                                                                                                                                                                                                                                         
wire [31:0]e42;                                                                                                                                                                                                                                         
wire [31:0]f42;                                                                                                                                                                                                                                         
wire [31:0]g42;
wire [31:0]h42;                                                                                                                                                                                                                                         
SHA256Node node42(a41,b41,c41,d41,e41,f41,g41,h41,a42,b42,c42,d42,e42,f42,g42,h42,k42,w42);                                                                                                                                                                     
wire [31:0]a43;                                                                                                                                                                                                                                         
wire [31:0]b43;                                                                                                                                                                                                                                         
wire [31:0]c43;                                                                                                                                                                                                                                         
wire [31:0]d43;                                                                                                                                                                                                                                         
wire [31:0]e43;                                                                                                                                                                                                                                         
wire [31:0]f43;                                                                                                                                                                                                                                         
wire [31:0]g43;
wire [31:0]h43;                                                                                                                                                                                                                                         
SHA256Node node43(a42,b42,c42,d42,e42,f42,g42,h42,a43,b43,c43,d43,e43,f43,g43,h43,k43,w43);                                                                                                                                                                     
wire [31:0]a44;                                                                                                                                                                                                                                         
wire [31:0]b44;                                                                                                                                                                                                                                         
wire [31:0]c44;                                                                                                                                                                                                                                         
wire [31:0]d44;                                                                                                                                                                                                                                         
wire [31:0]e44;                                                                                                                                                                                                                                         
wire [31:0]f44;                                                                                                                                                                                                                                         
wire [31:0]g44;
wire [31:0]h44;                                                                                                                                                                                                                                         
SHA256Node node44(a43,b43,c43,d43,e43,f43,g43,h43,a44,b44,c44,d44,e44,f44,g44,h44,k44,w44);
wire [31:0]a45;                                                                                                                                                                                                                                         
wire [31:0]b45;                                                                                                                                                                                                                                         
wire [31:0]c45;                                                                                                                                                                                                                                         
wire [31:0]d45;                                                                                                                                                                                                                                         
wire [31:0]e45;                                                                                                                                                                                                                                         
wire [31:0]f45;                                                                                                                                                                                                                                         
wire [31:0]g45;
wire [31:0]h45;                                                                                                                                                                                                                                         
SHA256Node node45(a44,b44,c44,d44,e44,f44,g44,h44,a45,b45,c45,d45,e45,f45,g45,h45,k45,w45);                                                                                                                                                                     
wire [31:0]a46;                                                                                                                                                                                                                                         
wire [31:0]b46;                                                                                                                                                                                                                                         
wire [31:0]c46;                                                                                                                                                                                                                                         
wire [31:0]d46;                                                                                                                                                                                                                                         
wire [31:0]e46;                                                                                                                                                                                                                                         
wire [31:0]f46;                                                                                                                                                                                                                                         
wire [31:0]g46;
wire [31:0]h46;                                                                                                                                                                                                                                         
SHA256Node node46(a45,b45,c45,d45,e45,f45,g45,h45,a46,b46,c46,d46,e46,f46,g46,h46,k46,w46);                                                                                                                                                                     
wire [31:0]a47;                                                                                                                                                                                                                                         
wire [31:0]b47;                                                                                                                                                                                                                                         
wire [31:0]c47;                                                                                                                                                                                                                                         
wire [31:0]d47;                                                                                                                                                                                                                                         
wire [31:0]e47;                                                                                                                                                                                                                                         
wire [31:0]f47;                                                                                                                                                                                                                                         
wire [31:0]g47;
wire [31:0]h47;                                                                                                                                                                                                                                         
SHA256Node node47(a46,b46,c46,d46,e46,f46,g46,h46,a47,b47,c47,d47,e47,f47,g47,h47,k47,w47);                                                                                                                                                                     
wire [31:0]a48;                                                                                                                                                                                                                                         
wire [31:0]b48;                                                                                                                                                                                                                                         
wire [31:0]c48;                                                                                                                                                                                                                                         
wire [31:0]d48;                                                                                                                                                                                                                                         
wire [31:0]e48;                                                                                                                                                                                                                                         
wire [31:0]f48;                                                                                                                                                                                                                                         
wire [31:0]g48;
wire [31:0]h48;                                                                                                                                                                                                                                         
SHA256Node node48(a47,b47,c47,d47,e47,f47,g47,h47,a48,b48,c48,d48,e48,f48,g48,h48,k48,w48);                                                                                                                                                                     
wire [31:0]a49;                                                                                                                                                                                                                                         
wire [31:0]b49;                                                                                                                                                                                                                                         
wire [31:0]c49;                                                                                                                                                                                                                                         
wire [31:0]d49;                                                                                                                                                                                                                                         
wire [31:0]e49;                                                                                                                                                                                                                                         
wire [31:0]f49;                                                                                                                                                                                                                                         
wire [31:0]g49;
wire [31:0]h49;                                                                                                                                                                                                                                         
SHA256Node node49(a48,b48,c48,d48,e48,f48,g48,h48,a49,b49,c49,d49,e49,f49,g49,h49,k49,w49);
wire [31:0]a50;                                                                                                                                                                                                                                         
wire [31:0]b50;                                                                                                                                                                                                                                         
wire [31:0]c50;                                                                                                                                                                                                                                         
wire [31:0]d50;                                                                                                                                                                                                                                         
wire [31:0]e50;                                                                                                                                                                                                                                         
wire [31:0]f50;                                                                                                                                                                                                                                         
wire [31:0]g50;
wire [31:0]h50;                                                                                                                                                                                                                                         
SHA256Node node50(a49,b49,c49,d49,e49,f49,g49,h49,a50,b50,c50,d50,e50,f50,g50,h50,k50,w50);                                                                                                                                                                     
wire [31:0]a51;                                                                                                                                                                                                                                         
wire [31:0]b51;                                                                                                                                                                                                                                         
wire [31:0]c51;                                                                                                                                                                                                                                         
wire [31:0]d51;                                                                                                                                                                                                                                         
wire [31:0]e51;                                                                                                                                                                                                                                         
wire [31:0]f51;                                                                                                                                                                                                                                         
wire [31:0]g51;
wire [31:0]h51;                                                                                                                                                                                                                                         
SHA256Node node51(a50,b50,c50,d50,e50,f50,g50,h50,a51,b51,c51,d51,e51,f51,g51,h51,k51,w51);                                                                                                                                                                     
wire [31:0]a52;                                                                                                                                                                                                                                         
wire [31:0]b52;                                                                                                                                                                                                                                         
wire [31:0]c52;                                                                                                                                                                                                                                         
wire [31:0]d52;                                                                                                                                                                                                                                         
wire [31:0]e52;                                                                                                                                                                                                                                         
wire [31:0]f52;                                                                                                                                                                                                                                         
wire [31:0]g52;
wire [31:0]h52;                                                                                                                                                                                                                                         
SHA256Node node52(a51,b51,c51,d51,e51,f51,g51,h51,a52,b52,c52,d52,e52,f52,g52,h52,k52,w52);                                                                                                                                                                     
wire [31:0]a53;                                                                                                                                                                                                                                         
wire [31:0]b53;                                                                                                                                                                                                                                         
wire [31:0]c53;                                                                                                                                                                                                                                         
wire [31:0]d53;                                                                                                                                                                                                                                         
wire [31:0]e53;                                                                                                                                                                                                                                         
wire [31:0]f53;                                                                                                                                                                                                                                         
wire [31:0]g53;
wire [31:0]h53;                                                                                                                                                                                                                                         
SHA256Node node53(a52,b52,c52,d52,e52,f52,g52,h52,a53,b53,c53,d53,e53,f53,g53,h53,k53,w53);                                                                                                                                                                     
wire [31:0]a54;                                                                                                                                                                                                                                         
wire [31:0]b54;                                                                                                                                                                                                                                         
wire [31:0]c54;                                                                                                                                                                                                                                         
wire [31:0]d54;                                                                                                                                                                                                                                         
wire [31:0]e54;                                                                                                                                                                                                                                         
wire [31:0]f54;                                                                                                                                                                                                                                         
wire [31:0]g54;
wire [31:0]h54;                                                                                                                                                                                                                                         
SHA256Node node54(a53,b53,c53,d53,e53,f53,g53,h53,a54,b54,c54,d54,e54,f54,g54,h54,k54,w54);
wire [31:0]a55;                                                                                                                                                                                                                                         
wire [31:0]b55;                                                                                                                                                                                                                                         
wire [31:0]c55;                                                                                                                                                                                                                                         
wire [31:0]d55;                                                                                                                                                                                                                                         
wire [31:0]e55;                                                                                                                                                                                                                                         
wire [31:0]f55;                                                                                                                                                                                                                                         
wire [31:0]g55;
wire [31:0]h55;                                                                                                                                                                                                                                         
SHA256Node node55(a54,b54,c54,d54,e54,f54,g54,h54,a55,b55,c55,d55,e55,f55,g55,h55,k55,w55);                                                                                                                                                                     
wire [31:0]a56;                                                                                                                                                                                                                                         
wire [31:0]b56;                                                                                                                                                                                                                                         
wire [31:0]c56;                                                                                                                                                                                                                                         
wire [31:0]d56;                                                                                                                                                                                                                                         
wire [31:0]e56;                                                                                                                                                                                                                                         
wire [31:0]f56;                                                                                                                                                                                                                                         
wire [31:0]g56;
wire [31:0]h56;                                                                                                                                                                                                                                         
SHA256Node node56(a55,b55,c55,d55,e55,f55,g55,h55,a56,b56,c56,d56,e56,f56,g56,h56,k56,w56);                                                                                                                                                                     
wire [31:0]a57;                                                                                                                                                                                                                                         
wire [31:0]b57;                                                                                                                                                                                                                                         
wire [31:0]c57;                                                                                                                                                                                                                                         
wire [31:0]d57;                                                                                                                                                                                                                                         
wire [31:0]e57;                                                                                                                                                                                                                                         
wire [31:0]f57;                                                                                                                                                                                                                                         
wire [31:0]g57;
wire [31:0]h57;                                                                                                                                                                                                                                         
SHA256Node node57(a56,b56,c56,d56,e56,f56,g56,h56,a57,b57,c57,d57,e57,f57,g57,h57,k57,w57);                                                                                                                                                                     
wire [31:0]a58;                                                                                                                                                                                                                                         
wire [31:0]b58;                                                                                                                                                                                                                                         
wire [31:0]c58;                                                                                                                                                                                                                                         
wire [31:0]d58;                                                                                                                                                                                                                                         
wire [31:0]e58;                                                                                                                                                                                                                                         
wire [31:0]f58;                                                                                                                                                                                                                                         
wire [31:0]g58;
wire [31:0]h58;                                                                                                                                                                                                                                         
SHA256Node node58(a57,b57,c57,d57,e57,f57,g57,h57,a58,b58,c58,d58,e58,f58,g58,h58,k58,w58);                                                                                                                                                                     
wire [31:0]a59;                                                                                                                                                                                                                                         
wire [31:0]b59;                                                                                                                                                                                                                                         
wire [31:0]c59;                                                                                                                                                                                                                                         
wire [31:0]d59;                                                                                                                                                                                                                                         
wire [31:0]e59;                                                                                                                                                                                                                                         
wire [31:0]f59;                                                                                                                                                                                                                                         
wire [31:0]g59;
wire [31:0]h59;                                                                                                                                                                                                                                         
SHA256Node node59(a58,b58,c58,d58,e58,f58,g58,h58,a59,b59,c59,d59,e59,f59,g59,h59,k59,w59);
wire [31:0]a60;                                                                                                                                                                                                                                         
wire [31:0]b60;                                                                                                                                                                                                                                         
wire [31:0]c60;                                                                                                                                                                                                                                         
wire [31:0]d60;                                                                                                                                                                                                                                         
wire [31:0]e60;                                                                                                                                                                                                                                         
wire [31:0]f60;                                                                                                                                                                                                                                         
wire [31:0]g60;
wire [31:0]h60;                                                                                                                                                                                                                                         
SHA256Node node60(a59,b59,c59,d59,e59,f59,g59,h59,a60,b60,c60,d60,e60,f60,g60,h60,k60,w60);                                                                                                                                                                     
wire [31:0]a61;                                                                                                                                                                                                                                         
wire [31:0]b61;                                                                                                                                                                                                                                         
wire [31:0]c61;                                                                                                                                                                                                                                         
wire [31:0]d61;                                                                                                                                                                                                                                         
wire [31:0]e61;                                                                                                                                                                                                                                         
wire [31:0]f61;                                                                                                                                                                                                                                         
wire [31:0]g61;
wire [31:0]h61;                                                                                                                                                                                                                                         
SHA256Node node61(a60,b60,c60,d60,e60,f60,g60,h60,a61,b61,c61,d61,e61,f61,g61,h61,k61,w61);                                                                                                                                                                     
wire [31:0]a62;                                                                                                                                                                                                                                         
wire [31:0]b62;                                                                                                                                                                                                                                         
wire [31:0]c62;                                                                                                                                                                                                                                         
wire [31:0]d62;                                                                                                                                                                                                                                         
wire [31:0]e62;                                                                                                                                                                                                                                         
wire [31:0]f62;                                                                                                                                                                                                                                         
wire [31:0]g62;
wire [31:0]h62;                                                                                                                                                                                                                                         
SHA256Node node62(a61,b61,c61,d61,e61,f61,g61,h61,a62,b62,c62,d62,e62,f62,g62,h62,k62,w62);                                                                                                                                                                     
wire [31:0]a63;                                                                                                                                                                                                                                         
wire [31:0]b63;                                                                                                                                                                                                                                         
wire [31:0]c63;                                                                                                                                                                                                                                         
wire [31:0]d63;                                                                                                                                                                                                                                         
wire [31:0]e63;                                                                                                                                                                                                                                         
wire [31:0]f63;                                                                                                                                                                                                                                         
wire [31:0]g63;
wire [31:0]h63;                                                                                                                                                                                                                                         
SHA256Node node63(a62,b62,c62,d62,e62,f62,g62,h62,a63,b63,c63,d63,e63,f63,g63,h63,k63,w63);                                                                                                                                                                                                                                                                                                                                                                                                              
SHA256Node node64(a63,b63,c63,d63,e63,f63,g63,h63,aout,bout,cout,dout,eout,fout,gout,hout,k64,w64);
//post nodes
wire [31:0]afinal;                                                                                                                                                                                                                                         
wire [31:0]bfinal;                                                                                                                                                                                                                                         
wire [31:0]cfinal;                                                                                                                                                                                                                                         
wire [31:0]dfinal;                                                                                                                                                                                                                                         
wire [31:0]efinal;                                                                                                                                                                                                                                         
wire [31:0]ffinal;                                                                                                                                                                                                                                         
wire [31:0]gfinal;
wire [31:0]hfinal;
assign afinal=aout+ainit;
assign bfinal=bout+binit;
assign cfinal=cout+cinit;
assign dfinal=dout+dinit;
assign efinal=eout+einit;
assign ffinal=fout+finit;
assign gfinal=gout+ginit;
assign hfinal=hout+hinit;
// final 256 bit output
assign out ={afinal,bfinal,cfinal,dfinal,efinal,ffinal,gfinal,hfinal};
endmodule
